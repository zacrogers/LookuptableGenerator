library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity sin_lut is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	addr     : in  std_logic_vector(23 downto 0);
	sin_out  : out std_logic_vector(23 downto 0)
);

end entity;


architecture rtl of sin_lut is

type rom_type is array (0 to 4096) of std_logic_vector (23  downto 0);

constant sin_ROM : rom_type :=
(
X"000000",X"003243",X"006487",X"0096cb",X"00c90f",X"00fb53",X"012d96",
X"015fda",X"01921d",X"01c45f",X"01f6a2",X"0228e4",X"025b26",X"028d68",
X"02bfa9",X"02f1ea",X"03242a",X"03566a",X"0388a9",X"03bae8",X"03ed26",
X"041f64",X"0451a1",X"0483dd",X"04b619",X"04e854",X"051a8e",X"054cc7",
X"057f00",X"05b137",X"05e36e",X"0615a4",X"0647d9",X"067a0d",X"06ac40",
X"06de72",X"0710a3",X"0742d3",X"077501",X"07a72f",X"07d95b",X"080b86",
X"083db0",X"086fd9",X"08a200",X"08d426",X"09064b",X"09386e",X"096a90",
X"099cb0",X"09cecf",X"0a00ec",X"0a3308",X"0a6522",X"0a973b",X"0ac952",
X"0afb68",X"0b2d7b",X"0b5f8d",X"0b919d",X"0bc3ac",X"0bf5b8",X"0c27c3",
X"0c59cc",X"0c8bd3",X"0cbdd8",X"0cefdb",X"0d21dc",X"0d53db",X"0d85d8",
X"0db7d3",X"0de9cc",X"0e1bc2",X"0e4db7",X"0e7fa9",X"0eb199",X"0ee387",
X"0f1572",X"0f475b",X"0f7942",X"0fab27",X"0fdd09",X"100ee8",X"1040c5",
X"1072a0",X"10a478",X"10d64d",X"110820",X"1139f0",X"116bbe",X"119d89",
X"11cf51",X"120116",X"1232d9",X"126499",X"129656",X"12c810",X"12f9c7",
X"132b7b",X"135d2d",X"138edb",X"13c087",X"13f22f",X"1423d4",X"145576",
X"148715",X"14b8b1",X"14ea4a",X"151bdf",X"154d71",X"157f00",X"15b08c",
X"15e214",X"161399",X"16451a",X"167698",X"16a813",X"16d98a",X"170afd",
X"173c6d",X"176dd9",X"179f42",X"17d0a7",X"180209",X"183366",X"1864c0",
X"189617",X"18c769",X"18f8b8",X"192a03",X"195b49",X"198c8c",X"19bdcb",
X"19ef07",X"1a203e",X"1a5171",X"1a82a0",X"1ab3cb",X"1ae4f1",X"1b1614",
X"1b4732",X"1b784d",X"1ba963",X"1bda74",X"1c0b82",X"1c3c8b",X"1c6d90",
X"1c9e90",X"1ccf8c",X"1d0084",X"1d3177",X"1d6265",X"1d934f",X"1dc435",
X"1df516",X"1e25f2",X"1e56ca",X"1e879d",X"1eb86b",X"1ee934",X"1f19f9",
X"1f4ab9",X"1f7b74",X"1fac2a",X"1fdcdc",X"200d88",X"203e30",X"206ed2",
X"209f70",X"20d008",X"21009c",X"21312a",X"2161b3",X"219237",X"21c2b6",
X"21f330",X"2223a4",X"225413",X"22847d",X"22b4e2",X"22e541",X"23159b",
X"2345ef",X"23763e",X"23a688",X"23d6cc",X"24070b",X"243743",X"246777",
X"2497a5",X"24c7cd",X"24f7ef",X"25280c",X"255823",X"258834",X"25b840",
X"25e845",X"261845",X"26483f",X"267833",X"26a821",X"26d809",X"2707eb",
X"2737c7",X"27679d",X"27976d",X"27c737",X"27f6fb",X"2826b9",X"285670",
X"288621",X"28b5cc",X"28e571",X"29150f",X"2944a7",X"297439",X"29a3c4",
X"29d349",X"2a02c7",X"2a323f",X"2a61b1",X"2a911b",X"2ac080",X"2aefdd",
X"2b1f34",X"2b4e85",X"2b7dcf",X"2bad12",X"2bdc4e",X"2c0b83",X"2c3ab2",
X"2c69da",X"2c98fb",X"2cc815",X"2cf729",X"2d2635",X"2d553a",X"2d8439",
X"2db330",X"2de221",X"2e110a",X"2e3fec",X"2e6ec7",X"2e9d9b",X"2ecc68",
X"2efb2d",X"2f29eb",X"2f58a2",X"2f8752",X"2fb5fa",X"2fe49b",X"301335",
X"3041c7",X"307052",X"309ed5",X"30cd51",X"30fbc5",X"312a31",X"315897",
X"3186f4",X"31b54a",X"31e398",X"3211df",X"32401d",X"326e54",X"329c84",
X"32caab",X"32f8cb",X"3326e2",X"3354f2",X"3382fa",X"33b0fa",X"33def2",
X"340ce2",X"343aca",X"3468aa",X"349682",X"34c452",X"34f219",X"351fd9",
X"354d90",X"357b3f",X"35a8e6",X"35d684",X"36041a",X"3631a8",X"365f2e",
X"368cab",X"36ba20",X"36e78c",X"3714f0",X"37424b",X"376f9e",X"379ce8",
X"37ca2a",X"37f763",X"382493",X"3851bb",X"387eda",X"38abf0",X"38d8fe",
X"390603",X"3932ff",X"395ff2",X"398cdd",X"39b9be",X"39e697",X"3a1367",
X"3a402d",X"3a6ceb",X"3a99a0",X"3ac64c",X"3af2ee",X"3b1f88",X"3b4c18",
X"3b78a0",X"3ba51e",X"3bd193",X"3bfdfe",X"3c2a61",X"3c56ba",X"3c830a",
X"3caf50",X"3cdb8e",X"3d07c1",X"3d33ec",X"3d600d",X"3d8c24",X"3db832",
X"3de437",X"3e1032",X"3e3c23",X"3e680b",X"3e93e9",X"3ebfbd",X"3eeb88",
X"3f1749",X"3f4301",X"3f6eae",X"3f9a52",X"3fc5ec",X"3ff17c",X"401d03",
X"40487f",X"4073f2",X"409f5a",X"40cab9",X"40f60d",X"412158",X"414c99",
X"4177cf",X"41a2fc",X"41ce1e",X"41f936",X"422444",X"424f48",X"427a41",
X"42a531",X"42d016",X"42faf0",X"4325c1",X"435087",X"437b42",X"43a5f4",
X"43d09a",X"43fb37",X"4425c9",X"445050",X"447acd",X"44a53f",X"44cfa7",
X"44fa04",X"452456",X"454e9e",X"4578db",X"45a30d",X"45cd35",X"45f752",
X"462164",X"464b6b",X"467568",X"469f59",X"46c940",X"46f31c",X"471cec",
X"4746b2",X"47706d",X"479a1d",X"47c3c2",X"47ed5b",X"4816ea",X"48406e",
X"4869e6",X"489353",X"48bcb5",X"48e60c",X"490f57",X"493898",X"4961cd",
X"498af6",X"49b415",X"49dd28",X"4a062f",X"4a2f2b",X"4a581c",X"4a8101",
X"4aa9db",X"4ad2a9",X"4afb6c",X"4b2423",X"4b4ccf",X"4b756f",X"4b9e03",
X"4bc68c",X"4bef09",X"4c177a",X"4c3fdf",X"4c6839",X"4c9087",X"4cb8c9",
X"4ce100",X"4d092a",X"4d3149",X"4d595b",X"4d8162",X"4da95d",X"4dd14c",
X"4df92f",X"4e2106",X"4e48d0",X"4e708f",X"4e9842",X"4ebfe8",X"4ee782",
X"4f0f11",X"4f3693",X"4f5e08",X"4f8572",X"4faccf",X"4fd420",X"4ffb65",
X"50229d",X"5049c9",X"5070e9",X"5097fc",X"50bf03",X"50e5fd",X"510ceb",
X"5133cc",X"515aa1",X"518169",X"51a825",X"51ced4",X"51f576",X"521c0c",
X"524295",X"526912",X"528f82",X"52b5e5",X"52dc3b",X"530285",X"5328c1",
X"534ef1",X"537514",X"539b2a",X"53c134",X"53e730",X"540d20",X"543302",
X"5458d7",X"547ea0",X"54a45b",X"54ca0a",X"54efab",X"55153f",X"553ac6",
X"556040",X"5585ad",X"55ab0d",X"55d05f",X"55f5a4",X"561adc",X"564007",
X"566524",X"568a34",X"56af37",X"56d42c",X"56f914",X"571dee",X"5742bc",
X"57677b",X"578c2d",X"57b0d2",X"57d569",X"57f9f2",X"581e6e",X"5842dd",
X"58673e",X"588b91",X"58afd6",X"58d40e",X"58f838",X"591c55",X"594063",
X"596464",X"598857",X"59ac3c",X"59d014",X"59f3de",X"5a1799",X"5a3b47",
X"5a5ee7",X"5a8279",X"5aa5fd",X"5ac973",X"5aecdb",X"5b1035",X"5b3381",
X"5b56bf",X"5b79ef",X"5b9d11",X"5bc024",X"5be32a",X"5c0621",X"5c290a",
X"5c4be5",X"5c6eb2",X"5c9170",X"5cb420",X"5cd6c2",X"5cf956",X"5d1bdb",
X"5d3e52",X"5d60ba",X"5d8314",X"5da560",X"5dc79d",X"5de9cc",X"5e0bec",
X"5e2dfe",X"5e5001",X"5e71f6",X"5e93dc",X"5eb5b3",X"5ed77c",X"5ef936",
X"5f1ae2",X"5f3c7f",X"5f5e0d",X"5f7f8d",X"5fa0fe",X"5fc260",X"5fe3b3",
X"6004f8",X"60262d",X"604754",X"60686c",X"608976",X"60aa70",X"60cb5b",
X"60ec38",X"610d05",X"612dc4",X"614e73",X"616f14",X"618fa5",X"61b028",
X"61d09b",X"61f100",X"621155",X"62319b",X"6251d2",X"6271fa",X"629213",
X"62b21c",X"62d216",X"62f201",X"6311dd",X"6331a9",X"635166",X"637114",
X"6390b3",X"63b042",X"63cfc2",X"63ef32",X"640e93",X"642de5",X"644d27",
X"646c59",X"648b7c",X"64aa90",X"64c994",X"64e889",X"65076e",X"652643",
X"654509",X"6563bf",X"658266",X"65a0fd",X"65bf84",X"65ddfb",X"65fc63",
X"661abb",X"663904",X"66573c",X"667565",X"66937e",X"66b187",X"66cf81",
X"66ed6a",X"670b44",X"67290e",X"6746c7",X"676471",X"67820b",X"679f95",
X"67bd0f",X"67da79",X"67f7d3",X"68151d",X"683257",X"684f81",X"686c9b",
X"6889a4",X"68a69e",X"68c387",X"68e061",X"68fd2a",X"6919e3",X"69368b",
X"695324",X"696fac",X"698c24",X"69a88c",X"69c4e3",X"69e12a",X"69fd61",
X"6a1987",X"6a359d",X"6a51a3",X"6a6d98",X"6a897d",X"6aa551",X"6ac115",
X"6adcc9",X"6af86c",X"6b13fe",X"6b2f80",X"6b4af2",X"6b6653",X"6b81a3",
X"6b9ce3",X"6bb812",X"6bd331",X"6bee3f",X"6c093c",X"6c2429",X"6c3f05",
X"6c59d0",X"6c748b",X"6c8f35",X"6ca9ce",X"6cc456",X"6cdece",X"6cf934",
X"6d138a",X"6d2dd0",X"6d4804",X"6d6227",X"6d7c3a",X"6d963c",X"6db02d",
X"6dca0d",X"6de3dc",X"6dfd9a",X"6e1747",X"6e30e3",X"6e4a6e",X"6e63e8",
X"6e7d51",X"6e96a9",X"6eaff0",X"6ec926",X"6ee24b",X"6efb5f",X"6f1461",
X"6f2d53",X"6f4633",X"6f5f02",X"6f77c0",X"6f906d",X"6fa909",X"6fc193",
X"6fda0c",X"6ff274",X"700acb",X"702310",X"703b44",X"705367",X"706b78",
X"708378",X"709b67",X"70b345",X"70cb11",X"70e2cb",X"70fa74",X"71120c",
X"712993",X"714108",X"71586b",X"716fbd",X"7186fd",X"719e2c",X"71b54a",
X"71cc56",X"71e350",X"71fa39",X"721110",X"7227d6",X"723e8a",X"72552c",
X"726bbd",X"72823c",X"7298a9",X"72af05",X"72c54f",X"72db88",X"72f1ae",
X"7307c3",X"731dc7",X"7333b8",X"734998",X"735f66",X"737522",X"738acc",
X"73a065",X"73b5eb",X"73cb60",X"73e0c3",X"73f614",X"740b53",X"742081",
X"74359c",X"744aa6",X"745f9d",X"747483",X"748957",X"749e18",X"74b2c8",
X"74c766",X"74dbf1",X"74f06b",X"7504d3",X"751928",X"752d6c",X"75419d",
X"7555bd",X"7569ca",X"757dc5",X"7591ae",X"75a585",X"75b94a",X"75ccfd",
X"75e09d",X"75f42c",X"7607a8",X"761b12",X"762e69",X"7641af",X"7654e2",
X"766803",X"767b12",X"768e0e",X"76a0f8",X"76b3d0",X"76c696",X"76d949",
X"76ebea",X"76fe79",X"7710f5",X"77235f",X"7735b6",X"7747fb",X"775a2e",
X"776c4e",X"777e5c",X"779058",X"77a241",X"77b417",X"77c5dc",X"77d78d",
X"77e92c",X"77fab9",X"780c33",X"781d9b",X"782ef0",X"784033",X"785163",
X"786280",X"78738b",X"788484",X"789569",X"78a63d",X"78b6fd",X"78c7ab",
X"78d846",X"78e8cf",X"78f945",X"7909a9",X"7919f9",X"792a37",X"793a63",
X"794a7c",X"795a82",X"796a75",X"797a55",X"798a23",X"7999de",X"79a987",
X"79b91c",X"79c89f",X"79d80f",X"79e76c",X"79f6b7",X"7a05ee",X"7a1513",
X"7a2425",X"7a3324",X"7a4210",X"7a50ea",X"7a5fb0",X"7a6e64",X"7a7d05",
X"7a8b93",X"7a9a0e",X"7aa876",X"7ab6cb",X"7ac50d",X"7ad33d",X"7ae159",
X"7aef63",X"7afd59",X"7b0b3d",X"7b190d",X"7b26cb",X"7b3475",X"7b420d",
X"7b4f92",X"7b5d03",X"7b6a62",X"7b77ad",X"7b84e6",X"7b920b",X"7b9f1d",
X"7bac1d",X"7bb909",X"7bc5e2",X"7bd2a8",X"7bdf5b",X"7bebfb",X"7bf888",
X"7c0501",X"7c1168",X"7c1dbb",X"7c29fb",X"7c3629",X"7c4242",X"7c4e49",
X"7c5a3d",X"7c661d",X"7c71ea",X"7c7da5",X"7c894b",X"7c94df",X"7ca05f",
X"7cabcd",X"7cb727",X"7cc26d",X"7ccda1",X"7cd8c1",X"7ce3ce",X"7ceec8",
X"7cf9ae",X"7d0482",X"7d0f42",X"7d19ee",X"7d2488",X"7d2f0e",X"7d3980",
X"7d43e0",X"7d4e2c",X"7d5865",X"7d628a",X"7d6c9c",X"7d769b",X"7d8087",
X"7d8a5f",X"7d9423",X"7d9dd5",X"7da773",X"7db0fd",X"7dba75",X"7dc3d9",
X"7dcd29",X"7dd666",X"7ddf90",X"7de8a6",X"7df1a9",X"7dfa98",X"7e0374",
X"7e0c3d",X"7e14f2",X"7e1d93",X"7e2622",X"7e2e9c",X"7e3704",X"7e3f57",
X"7e4798",X"7e4fc5",X"7e57de",X"7e5fe4",X"7e67d7",X"7e6fb5",X"7e7781",
X"7e7f39",X"7e86dd",X"7e8e6e",X"7e95ec",X"7e9d55",X"7ea4ac",X"7eabef",
X"7eb31e",X"7eba3a",X"7ec142",X"7ec837",X"7ecf18",X"7ed5e5",X"7edc9f",
X"7ee346",X"7ee9d9",X"7ef058",X"7ef6c4",X"7efd1c",X"7f0360",X"7f0991",
X"7f0faf",X"7f15b8",X"7f1baf",X"7f2191",X"7f2760",X"7f2d1c",X"7f32c3",
X"7f3857",X"7f3dd8",X"7f4345",X"7f489e",X"7f4de4",X"7f5316",X"7f5834",
X"7f5d3f",X"7f6236",X"7f671a",X"7f6be9",X"7f70a5",X"7f754e",X"7f79e3",
X"7f7e64",X"7f82d2",X"7f872b",X"7f8b72",X"7f8fa4",X"7f93c3",X"7f97ce",
X"7f9bc6",X"7f9faa",X"7fa37a",X"7fa736",X"7faadf",X"7fae74",X"7fb1f5",
X"7fb563",X"7fb8bd",X"7fbc04",X"7fbf36",X"7fc255",X"7fc560",X"7fc858",
X"7fcb3c",X"7fce0c",X"7fd0c8",X"7fd371",X"7fd606",X"7fd887",X"7fdaf5",
X"7fdd4e",X"7fdf95",X"7fe1c7",X"7fe3e6",X"7fe5f1",X"7fe7e8",X"7fe9cb",
X"7feb9b",X"7fed57",X"7feeff",X"7ff094",X"7ff215",X"7ff382",X"7ff4db",
X"7ff621",X"7ff753",X"7ff871",X"7ff97c",X"7ffa72",X"7ffb55",X"7ffc25",
X"7ffce0",X"7ffd88",X"7ffe1c",X"7ffe9c",X"7fff09",X"7fff62",X"7fffa7",
X"7fffd8",X"7ffff6",X"800000",X"7ffff6",X"7fffd8",X"7fffa7",X"7fff62",
X"7fff09",X"7ffe9c",X"7ffe1c",X"7ffd88",X"7ffce0",X"7ffc25",X"7ffb55",
X"7ffa72",X"7ff97c",X"7ff871",X"7ff753",X"7ff621",X"7ff4db",X"7ff382",
X"7ff215",X"7ff094",X"7feeff",X"7fed57",X"7feb9b",X"7fe9cb",X"7fe7e8",
X"7fe5f1",X"7fe3e6",X"7fe1c7",X"7fdf95",X"7fdd4e",X"7fdaf5",X"7fd887",
X"7fd606",X"7fd371",X"7fd0c8",X"7fce0c",X"7fcb3c",X"7fc858",X"7fc560",
X"7fc255",X"7fbf36",X"7fbc04",X"7fb8bd",X"7fb563",X"7fb1f5",X"7fae74",
X"7faadf",X"7fa736",X"7fa37a",X"7f9faa",X"7f9bc6",X"7f97ce",X"7f93c3",
X"7f8fa4",X"7f8b72",X"7f872b",X"7f82d2",X"7f7e64",X"7f79e3",X"7f754e",
X"7f70a5",X"7f6be9",X"7f671a",X"7f6236",X"7f5d3f",X"7f5834",X"7f5316",
X"7f4de4",X"7f489e",X"7f4345",X"7f3dd8",X"7f3857",X"7f32c3",X"7f2d1c",
X"7f2760",X"7f2191",X"7f1baf",X"7f15b8",X"7f0faf",X"7f0991",X"7f0360",
X"7efd1c",X"7ef6c4",X"7ef058",X"7ee9d9",X"7ee346",X"7edc9f",X"7ed5e5",
X"7ecf18",X"7ec837",X"7ec142",X"7eba3a",X"7eb31e",X"7eabef",X"7ea4ac",
X"7e9d55",X"7e95ec",X"7e8e6e",X"7e86dd",X"7e7f39",X"7e7781",X"7e6fb5",
X"7e67d7",X"7e5fe4",X"7e57de",X"7e4fc5",X"7e4798",X"7e3f57",X"7e3704",
X"7e2e9c",X"7e2622",X"7e1d93",X"7e14f2",X"7e0c3d",X"7e0374",X"7dfa98",
X"7df1a9",X"7de8a6",X"7ddf90",X"7dd666",X"7dcd29",X"7dc3d9",X"7dba75",
X"7db0fd",X"7da773",X"7d9dd5",X"7d9423",X"7d8a5f",X"7d8087",X"7d769b",
X"7d6c9c",X"7d628a",X"7d5865",X"7d4e2c",X"7d43e0",X"7d3980",X"7d2f0e",
X"7d2488",X"7d19ee",X"7d0f42",X"7d0482",X"7cf9ae",X"7ceec8",X"7ce3ce",
X"7cd8c1",X"7ccda1",X"7cc26d",X"7cb727",X"7cabcd",X"7ca05f",X"7c94df",
X"7c894b",X"7c7da5",X"7c71ea",X"7c661d",X"7c5a3d",X"7c4e49",X"7c4242",
X"7c3629",X"7c29fb",X"7c1dbb",X"7c1168",X"7c0501",X"7bf888",X"7bebfb",
X"7bdf5b",X"7bd2a8",X"7bc5e2",X"7bb909",X"7bac1d",X"7b9f1d",X"7b920b",
X"7b84e6",X"7b77ad",X"7b6a62",X"7b5d03",X"7b4f92",X"7b420d",X"7b3475",
X"7b26cb",X"7b190d",X"7b0b3d",X"7afd59",X"7aef63",X"7ae159",X"7ad33d",
X"7ac50d",X"7ab6cb",X"7aa876",X"7a9a0e",X"7a8b93",X"7a7d05",X"7a6e64",
X"7a5fb0",X"7a50ea",X"7a4210",X"7a3324",X"7a2425",X"7a1513",X"7a05ee",
X"79f6b7",X"79e76c",X"79d80f",X"79c89f",X"79b91c",X"79a987",X"7999de",
X"798a23",X"797a55",X"796a75",X"795a82",X"794a7c",X"793a63",X"792a37",
X"7919f9",X"7909a9",X"78f945",X"78e8cf",X"78d846",X"78c7ab",X"78b6fd",
X"78a63d",X"789569",X"788484",X"78738b",X"786280",X"785163",X"784033",
X"782ef0",X"781d9b",X"780c33",X"77fab9",X"77e92c",X"77d78d",X"77c5dc",
X"77b417",X"77a241",X"779058",X"777e5c",X"776c4e",X"775a2e",X"7747fb",
X"7735b6",X"77235f",X"7710f5",X"76fe79",X"76ebea",X"76d949",X"76c696",
X"76b3d0",X"76a0f8",X"768e0e",X"767b12",X"766803",X"7654e2",X"7641af",
X"762e69",X"761b12",X"7607a8",X"75f42c",X"75e09d",X"75ccfd",X"75b94a",
X"75a585",X"7591ae",X"757dc5",X"7569ca",X"7555bd",X"75419d",X"752d6c",
X"751928",X"7504d3",X"74f06b",X"74dbf1",X"74c766",X"74b2c8",X"749e18",
X"748957",X"747483",X"745f9d",X"744aa6",X"74359c",X"742081",X"740b53",
X"73f614",X"73e0c3",X"73cb60",X"73b5eb",X"73a065",X"738acc",X"737522",
X"735f66",X"734998",X"7333b8",X"731dc7",X"7307c3",X"72f1ae",X"72db88",
X"72c54f",X"72af05",X"7298a9",X"72823c",X"726bbd",X"72552c",X"723e8a",
X"7227d6",X"721110",X"71fa39",X"71e350",X"71cc56",X"71b54a",X"719e2c",
X"7186fd",X"716fbd",X"71586b",X"714108",X"712993",X"71120c",X"70fa74",
X"70e2cb",X"70cb11",X"70b345",X"709b67",X"708378",X"706b78",X"705367",
X"703b44",X"702310",X"700acb",X"6ff274",X"6fda0c",X"6fc193",X"6fa909",
X"6f906d",X"6f77c0",X"6f5f02",X"6f4633",X"6f2d53",X"6f1461",X"6efb5f",
X"6ee24b",X"6ec926",X"6eaff0",X"6e96a9",X"6e7d51",X"6e63e8",X"6e4a6e",
X"6e30e3",X"6e1747",X"6dfd9a",X"6de3dc",X"6dca0d",X"6db02d",X"6d963c",
X"6d7c3a",X"6d6227",X"6d4804",X"6d2dd0",X"6d138a",X"6cf934",X"6cdece",
X"6cc456",X"6ca9ce",X"6c8f35",X"6c748b",X"6c59d0",X"6c3f05",X"6c2429",
X"6c093c",X"6bee3f",X"6bd331",X"6bb812",X"6b9ce3",X"6b81a3",X"6b6653",
X"6b4af2",X"6b2f80",X"6b13fe",X"6af86c",X"6adcc9",X"6ac115",X"6aa551",
X"6a897d",X"6a6d98",X"6a51a3",X"6a359d",X"6a1987",X"69fd61",X"69e12a",
X"69c4e3",X"69a88c",X"698c24",X"696fac",X"695324",X"69368b",X"6919e3",
X"68fd2a",X"68e061",X"68c387",X"68a69e",X"6889a4",X"686c9b",X"684f81",
X"683257",X"68151d",X"67f7d3",X"67da79",X"67bd0f",X"679f95",X"67820b",
X"676471",X"6746c7",X"67290e",X"670b44",X"66ed6a",X"66cf81",X"66b187",
X"66937e",X"667565",X"66573c",X"663904",X"661abb",X"65fc63",X"65ddfb",
X"65bf84",X"65a0fd",X"658266",X"6563bf",X"654509",X"652643",X"65076e",
X"64e889",X"64c994",X"64aa90",X"648b7c",X"646c59",X"644d27",X"642de5",
X"640e93",X"63ef32",X"63cfc2",X"63b042",X"6390b3",X"637114",X"635166",
X"6331a9",X"6311dd",X"62f201",X"62d216",X"62b21c",X"629213",X"6271fa",
X"6251d2",X"62319b",X"621155",X"61f100",X"61d09b",X"61b028",X"618fa5",
X"616f14",X"614e73",X"612dc4",X"610d05",X"60ec38",X"60cb5b",X"60aa70",
X"608976",X"60686c",X"604754",X"60262d",X"6004f8",X"5fe3b3",X"5fc260",
X"5fa0fe",X"5f7f8d",X"5f5e0d",X"5f3c7f",X"5f1ae2",X"5ef936",X"5ed77c",
X"5eb5b3",X"5e93dc",X"5e71f6",X"5e5001",X"5e2dfe",X"5e0bec",X"5de9cc",
X"5dc79d",X"5da560",X"5d8314",X"5d60ba",X"5d3e52",X"5d1bdb",X"5cf956",
X"5cd6c2",X"5cb420",X"5c9170",X"5c6eb2",X"5c4be5",X"5c290a",X"5c0621",
X"5be32a",X"5bc024",X"5b9d11",X"5b79ef",X"5b56bf",X"5b3381",X"5b1035",
X"5aecdb",X"5ac973",X"5aa5fd",X"5a8279",X"5a5ee7",X"5a3b47",X"5a1799",
X"59f3de",X"59d014",X"59ac3c",X"598857",X"596464",X"594063",X"591c55",
X"58f838",X"58d40e",X"58afd6",X"588b91",X"58673e",X"5842dd",X"581e6e",
X"57f9f2",X"57d569",X"57b0d2",X"578c2d",X"57677b",X"5742bc",X"571dee",
X"56f914",X"56d42c",X"56af37",X"568a34",X"566524",X"564007",X"561adc",
X"55f5a4",X"55d05f",X"55ab0d",X"5585ad",X"556040",X"553ac6",X"55153f",
X"54efab",X"54ca0a",X"54a45b",X"547ea0",X"5458d7",X"543302",X"540d20",
X"53e730",X"53c134",X"539b2a",X"537514",X"534ef1",X"5328c1",X"530285",
X"52dc3b",X"52b5e5",X"528f82",X"526912",X"524295",X"521c0c",X"51f576",
X"51ced4",X"51a825",X"518169",X"515aa1",X"5133cc",X"510ceb",X"50e5fd",
X"50bf03",X"5097fc",X"5070e9",X"5049c9",X"50229d",X"4ffb65",X"4fd420",
X"4faccf",X"4f8572",X"4f5e08",X"4f3693",X"4f0f11",X"4ee782",X"4ebfe8",
X"4e9842",X"4e708f",X"4e48d0",X"4e2106",X"4df92f",X"4dd14c",X"4da95d",
X"4d8162",X"4d595b",X"4d3149",X"4d092a",X"4ce100",X"4cb8c9",X"4c9087",
X"4c6839",X"4c3fdf",X"4c177a",X"4bef09",X"4bc68c",X"4b9e03",X"4b756f",
X"4b4ccf",X"4b2423",X"4afb6c",X"4ad2a9",X"4aa9db",X"4a8101",X"4a581c",
X"4a2f2b",X"4a062f",X"49dd28",X"49b415",X"498af6",X"4961cd",X"493898",
X"490f57",X"48e60c",X"48bcb5",X"489353",X"4869e6",X"48406e",X"4816ea",
X"47ed5b",X"47c3c2",X"479a1d",X"47706d",X"4746b2",X"471cec",X"46f31c",
X"46c940",X"469f59",X"467568",X"464b6b",X"462164",X"45f752",X"45cd35",
X"45a30d",X"4578db",X"454e9e",X"452456",X"44fa04",X"44cfa7",X"44a53f",
X"447acd",X"445050",X"4425c9",X"43fb37",X"43d09a",X"43a5f4",X"437b42",
X"435087",X"4325c1",X"42faf0",X"42d016",X"42a531",X"427a41",X"424f48",
X"422444",X"41f936",X"41ce1e",X"41a2fc",X"4177cf",X"414c99",X"412158",
X"40f60d",X"40cab9",X"409f5a",X"4073f2",X"40487f",X"401d03",X"3ff17c",
X"3fc5ec",X"3f9a52",X"3f6eae",X"3f4301",X"3f1749",X"3eeb88",X"3ebfbd",
X"3e93e9",X"3e680b",X"3e3c23",X"3e1032",X"3de437",X"3db832",X"3d8c24",
X"3d600d",X"3d33ec",X"3d07c1",X"3cdb8e",X"3caf50",X"3c830a",X"3c56ba",
X"3c2a61",X"3bfdfe",X"3bd193",X"3ba51e",X"3b78a0",X"3b4c18",X"3b1f88",
X"3af2ee",X"3ac64c",X"3a99a0",X"3a6ceb",X"3a402d",X"3a1367",X"39e697",
X"39b9be",X"398cdd",X"395ff2",X"3932ff",X"390603",X"38d8fe",X"38abf0",
X"387eda",X"3851bb",X"382493",X"37f763",X"37ca2a",X"379ce8",X"376f9e",
X"37424b",X"3714f0",X"36e78c",X"36ba20",X"368cab",X"365f2e",X"3631a8",
X"36041a",X"35d684",X"35a8e6",X"357b3f",X"354d90",X"351fd9",X"34f219",
X"34c452",X"349682",X"3468aa",X"343aca",X"340ce2",X"33def2",X"33b0fa",
X"3382fa",X"3354f2",X"3326e2",X"32f8cb",X"32caab",X"329c84",X"326e54",
X"32401d",X"3211df",X"31e398",X"31b54a",X"3186f4",X"315897",X"312a31",
X"30fbc5",X"30cd51",X"309ed5",X"307052",X"3041c7",X"301335",X"2fe49b",
X"2fb5fa",X"2f8752",X"2f58a2",X"2f29eb",X"2efb2d",X"2ecc68",X"2e9d9b",
X"2e6ec7",X"2e3fec",X"2e110a",X"2de221",X"2db330",X"2d8439",X"2d553a",
X"2d2635",X"2cf729",X"2cc815",X"2c98fb",X"2c69da",X"2c3ab2",X"2c0b83",
X"2bdc4e",X"2bad12",X"2b7dcf",X"2b4e85",X"2b1f34",X"2aefdd",X"2ac080",
X"2a911b",X"2a61b1",X"2a323f",X"2a02c7",X"29d349",X"29a3c4",X"297439",
X"2944a7",X"29150f",X"28e571",X"28b5cc",X"288621",X"285670",X"2826b9",
X"27f6fb",X"27c737",X"27976d",X"27679d",X"2737c7",X"2707eb",X"26d809",
X"26a821",X"267833",X"26483f",X"261845",X"25e845",X"25b840",X"258834",
X"255823",X"25280c",X"24f7ef",X"24c7cd",X"2497a5",X"246777",X"243743",
X"24070b",X"23d6cc",X"23a688",X"23763e",X"2345ef",X"23159b",X"22e541",
X"22b4e2",X"22847d",X"225413",X"2223a4",X"21f330",X"21c2b6",X"219237",
X"2161b3",X"21312a",X"21009c",X"20d008",X"209f70",X"206ed2",X"203e30",
X"200d88",X"1fdcdc",X"1fac2a",X"1f7b74",X"1f4ab9",X"1f19f9",X"1ee934",
X"1eb86b",X"1e879d",X"1e56ca",X"1e25f2",X"1df516",X"1dc435",X"1d934f",
X"1d6265",X"1d3177",X"1d0084",X"1ccf8c",X"1c9e90",X"1c6d90",X"1c3c8b",
X"1c0b82",X"1bda74",X"1ba963",X"1b784d",X"1b4732",X"1b1614",X"1ae4f1",
X"1ab3cb",X"1a82a0",X"1a5171",X"1a203e",X"19ef07",X"19bdcb",X"198c8c",
X"195b49",X"192a03",X"18f8b8",X"18c769",X"189617",X"1864c0",X"183366",
X"180209",X"17d0a7",X"179f42",X"176dd9",X"173c6d",X"170afd",X"16d98a",
X"16a813",X"167698",X"16451a",X"161399",X"15e214",X"15b08c",X"157f00",
X"154d71",X"151bdf",X"14ea4a",X"14b8b1",X"148715",X"145576",X"1423d4",
X"13f22f",X"13c087",X"138edb",X"135d2d",X"132b7b",X"12f9c7",X"12c810",
X"129656",X"126499",X"1232d9",X"120116",X"11cf51",X"119d89",X"116bbe",
X"1139f0",X"110820",X"10d64d",X"10a478",X"1072a0",X"1040c5",X"100ee8",
X"0fdd09",X"0fab27",X"0f7942",X"0f475b",X"0f1572",X"0ee387",X"0eb199",
X"0e7fa9",X"0e4db7",X"0e1bc2",X"0de9cc",X"0db7d3",X"0d85d8",X"0d53db",
X"0d21dc",X"0cefdb",X"0cbdd8",X"0c8bd3",X"0c59cc",X"0c27c3",X"0bf5b8",
X"0bc3ac",X"0b919d",X"0b5f8d",X"0b2d7b",X"0afb68",X"0ac952",X"0a973b",
X"0a6522",X"0a3308",X"0a00ec",X"09cecf",X"099cb0",X"096a90",X"09386e",
X"09064b",X"08d426",X"08a200",X"086fd9",X"083db0",X"080b86",X"07d95b",
X"07a72f",X"077501",X"0742d3",X"0710a3",X"06de72",X"06ac40",X"067a0d",
X"0647d9",X"0615a4",X"05e36e",X"05b137",X"057f00",X"054cc7",X"051a8e",
X"04e854",X"04b619",X"0483dd",X"0451a1",X"041f64",X"03ed26",X"03bae8",
X"0388a9",X"03566a",X"03242a",X"02f1ea",X"02bfa9",X"028d68",X"025b26",
X"0228e4",X"01f6a2",X"01c45f",X"01921d",X"015fda",X"012d96",X"00fb53",
X"00c90f",X"0096cb",X"006487",X"003243",X"000000",X"ffcdbd",X"ff9b79",
X"ff6935",X"ff36f1",X"ff04ad",X"fed26a",X"fea026",X"fe6de3",X"fe3ba1",
X"fe095e",X"fdd71c",X"fda4da",X"fd7298",X"fd4057",X"fd0e16",X"fcdbd6",
X"fca996",X"fc7757",X"fc4518",X"fc12da",X"fbe09c",X"fbae5f",X"fb7c23",
X"fb49e7",X"fb17ac",X"fae572",X"fab339",X"fa8100",X"fa4ec9",X"fa1c92",
X"f9ea5c",X"f9b827",X"f985f3",X"f953c0",X"f9218e",X"f8ef5d",X"f8bd2d",
X"f88aff",X"f858d1",X"f826a5",X"f7f47a",X"f7c250",X"f79027",X"f75e00",
X"f72bda",X"f6f9b5",X"f6c792",X"f69570",X"f66350",X"f63131",X"f5ff14",
X"f5ccf8",X"f59ade",X"f568c5",X"f536ae",X"f50498",X"f4d285",X"f4a073",
X"f46e63",X"f43c54",X"f40a48",X"f3d83d",X"f3a634",X"f3742d",X"f34228",
X"f31025",X"f2de24",X"f2ac25",X"f27a28",X"f2482d",X"f21634",X"f1e43e",
X"f1b249",X"f18057",X"f14e67",X"f11c79",X"f0ea8e",X"f0b8a5",X"f086be",
X"f054d9",X"f022f7",X"eff118",X"efbf3b",X"ef8d60",X"ef5b88",X"ef29b3",
X"eef7e0",X"eec610",X"ee9442",X"ee6277",X"ee30af",X"edfeea",X"edcd27",
X"ed9b67",X"ed69aa",X"ed37f0",X"ed0639",X"ecd485",X"eca2d3",X"ec7125",
X"ec3f79",X"ec0dd1",X"ebdc2c",X"ebaa8a",X"eb78eb",X"eb474f",X"eb15b6",
X"eae421",X"eab28f",X"ea8100",X"ea4f74",X"ea1dec",X"e9ec67",X"e9bae6",
X"e98968",X"e957ed",X"e92676",X"e8f503",X"e8c393",X"e89227",X"e860be",
X"e82f59",X"e7fdf7",X"e7cc9a",X"e79b40",X"e769e9",X"e73897",X"e70748",
X"e6d5fd",X"e6a4b7",X"e67374",X"e64235",X"e610f9",X"e5dfc2",X"e5ae8f",
X"e57d60",X"e54c35",X"e51b0f",X"e4e9ec",X"e4b8ce",X"e487b3",X"e4569d",
X"e4258c",X"e3f47e",X"e3c375",X"e39270",X"e36170",X"e33074",X"e2ff7c",
X"e2ce89",X"e29d9b",X"e26cb1",X"e23bcb",X"e20aea",X"e1da0e",X"e1a936",
X"e17863",X"e14795",X"e116cc",X"e0e607",X"e0b547",X"e0848c",X"e053d6",
X"e02324",X"dff278",X"dfc1d0",X"df912e",X"df6090",X"df2ff8",X"deff64",
X"deced6",X"de9e4d",X"de6dc9",X"de3d4a",X"de0cd0",X"dddc5c",X"ddabed",
X"dd7b83",X"dd4b1e",X"dd1abf",X"dcea65",X"dcba11",X"dc89c2",X"dc5978",
X"dc2934",X"dbf8f5",X"dbc8bd",X"db9889",X"db685b",X"db3833",X"db0811",
X"dad7f4",X"daa7dd",X"da77cc",X"da47c0",X"da17bb",X"d9e7bb",X"d9b7c1",
X"d987cd",X"d957df",X"d927f7",X"d8f815",X"d8c839",X"d89863",X"d86893",
X"d838c9",X"d80905",X"d7d947",X"d7a990",X"d779df",X"d74a34",X"d71a8f",
X"d6eaf1",X"d6bb59",X"d68bc7",X"d65c3c",X"d62cb7",X"d5fd39",X"d5cdc1",
X"d59e4f",X"d56ee5",X"d53f80",X"d51023",X"d4e0cc",X"d4b17b",X"d48231",
X"d452ee",X"d423b2",X"d3f47d",X"d3c54e",X"d39626",X"d36705",X"d337eb",
X"d308d7",X"d2d9cb",X"d2aac6",X"d27bc7",X"d24cd0",X"d21ddf",X"d1eef6",
X"d1c014",X"d19139",X"d16265",X"d13398",X"d104d3",X"d0d615",X"d0a75e",
X"d078ae",X"d04a06",X"d01b65",X"cfeccb",X"cfbe39",X"cf8fae",X"cf612b",
X"cf32af",X"cf043b",X"ced5cf",X"cea769",X"ce790c",X"ce4ab6",X"ce1c68",
X"cdee21",X"cdbfe3",X"cd91ac",X"cd637c",X"cd3555",X"cd0735",X"ccd91e",
X"ccab0e",X"cc7d06",X"cc4f06",X"cc210e",X"cbf31e",X"cbc536",X"cb9756",
X"cb697e",X"cb3bae",X"cb0de7",X"cae027",X"cab270",X"ca84c1",X"ca571a",
X"ca297c",X"c9fbe6",X"c9ce58",X"c9a0d2",X"c97355",X"c945e0",X"c91874",
X"c8eb10",X"c8bdb5",X"c89062",X"c86318",X"c835d6",X"c8089d",X"c7db6d",
X"c7ae45",X"c78126",X"c75410",X"c72702",X"c6f9fd",X"c6cd01",X"c6a00e",
X"c67323",X"c64642",X"c61969",X"c5ec99",X"c5bfd3",X"c59315",X"c56660",
X"c539b4",X"c50d12",X"c4e078",X"c4b3e8",X"c48760",X"c45ae2",X"c42e6d",
X"c40202",X"c3d59f",X"c3a946",X"c37cf6",X"c350b0",X"c32472",X"c2f83f",
X"c2cc14",X"c29ff3",X"c273dc",X"c247ce",X"c21bc9",X"c1efce",X"c1c3dd",
X"c197f5",X"c16c17",X"c14043",X"c11478",X"c0e8b7",X"c0bcff",X"c09152",
X"c065ae",X"c03a14",X"c00e84",X"bfe2fd",X"bfb781",X"bf8c0e",X"bf60a6",
X"bf3547",X"bf09f3",X"bedea8",X"beb367",X"be8831",X"be5d04",X"be31e2",
X"be06ca",X"bddbbc",X"bdb0b8",X"bd85bf",X"bd5acf",X"bd2fea",X"bd0510",
X"bcda3f",X"bcaf79",X"bc84be",X"bc5a0c",X"bc2f66",X"bc04c9",X"bbda37",
X"bbafb0",X"bb8533",X"bb5ac1",X"bb3059",X"bb05fc",X"badbaa",X"bab162",
X"ba8725",X"ba5cf3",X"ba32cb",X"ba08ae",X"b9de9c",X"b9b495",X"b98a98",
X"b960a7",X"b936c0",X"b90ce4",X"b8e314",X"b8b94e",X"b88f93",X"b865e3",
X"b83c3e",X"b812a5",X"b7e916",X"b7bf92",X"b7961a",X"b76cad",X"b7434b",
X"b719f4",X"b6f0a9",X"b6c768",X"b69e33",X"b6750a",X"b64beb",X"b622d8",
X"b5f9d1",X"b5d0d5",X"b5a7e4",X"b57eff",X"b55625",X"b52d57",X"b50494",
X"b4dbdd",X"b4b331",X"b48a91",X"b461fd",X"b43974",X"b410f7",X"b3e886",
X"b3c021",X"b397c7",X"b36f79",X"b34737",X"b31f00",X"b2f6d6",X"b2ceb7",
X"b2a6a5",X"b27e9e",X"b256a3",X"b22eb4",X"b206d1",X"b1defa",X"b1b730",
X"b18f71",X"b167be",X"b14018",X"b1187e",X"b0f0ef",X"b0c96d",X"b0a1f8",
X"b07a8e",X"b05331",X"b02be0",X"b0049b",X"afdd63",X"afb637",X"af8f17",
X"af6804",X"af40fd",X"af1a03",X"aef315",X"aecc34",X"aea55f",X"ae7e97",
X"ae57db",X"ae312c",X"ae0a8a",X"ade3f4",X"adbd6b",X"ad96ee",X"ad707e",
X"ad4a1b",X"ad23c5",X"acfd7b",X"acd73f",X"acb10f",X"ac8aec",X"ac64d6",
X"ac3ecc",X"ac18d0",X"abf2e0",X"abccfe",X"aba729",X"ab8160",X"ab5ba5",
X"ab35f6",X"ab1055",X"aaeac1",X"aac53a",X"aa9fc0",X"aa7a53",X"aa54f3",
X"aa2fa1",X"aa0a5c",X"a9e524",X"a9bff9",X"a99adc",X"a975cc",X"a950c9",
X"a92bd4",X"a906ec",X"a8e212",X"a8bd44",X"a89885",X"a873d3",X"a84f2e",
X"a82a97",X"a8060e",X"a7e192",X"a7bd23",X"a798c2",X"a7746f",X"a7502a",
X"a72bf2",X"a707c8",X"a6e3ab",X"a6bf9d",X"a69b9c",X"a677a9",X"a653c4",
X"a62fec",X"a60c22",X"a5e867",X"a5c4b9",X"a5a119",X"a57d87",X"a55a03",
X"a5368d",X"a51325",X"a4efcb",X"a4cc7f",X"a4a941",X"a48611",X"a462ef",
X"a43fdc",X"a41cd6",X"a3f9df",X"a3d6f6",X"a3b41b",X"a3914e",X"a36e90",
X"a34be0",X"a3293e",X"a306aa",X"a2e425",X"a2c1ae",X"a29f46",X"a27cec",
X"a25aa0",X"a23863",X"a21634",X"a1f414",X"a1d202",X"a1afff",X"a18e0a",
X"a16c24",X"a14a4d",X"a12884",X"a106ca",X"a0e51e",X"a0c381",X"a0a1f3",
X"a08073",X"a05f02",X"a03da0",X"a01c4d",X"9ffb08",X"9fd9d3",X"9fb8ac",
X"9f9794",X"9f768a",X"9f5590",X"9f34a5",X"9f13c8",X"9ef2fb",X"9ed23c",
X"9eb18d",X"9e90ec",X"9e705b",X"9e4fd8",X"9e2f65",X"9e0f00",X"9deeab",
X"9dce65",X"9dae2e",X"9d8e06",X"9d6ded",X"9d4de4",X"9d2dea",X"9d0dff",
X"9cee23",X"9cce57",X"9cae9a",X"9c8eec",X"9c6f4d",X"9c4fbe",X"9c303e",
X"9c10ce",X"9bf16d",X"9bd21b",X"9bb2d9",X"9b93a7",X"9b7484",X"9b5570",
X"9b366c",X"9b1777",X"9af892",X"9ad9bd",X"9abaf7",X"9a9c41",X"9a7d9a",
X"9a5f03",X"9a407c",X"9a2205",X"9a039d",X"99e545",X"99c6fc",X"99a8c4",
X"998a9b",X"996c82",X"994e79",X"99307f",X"991296",X"98f4bc",X"98d6f2",
X"98b939",X"989b8f",X"987df5",X"98606b",X"9842f1",X"982587",X"98082d",
X"97eae3",X"97cda9",X"97b07f",X"979365",X"97765c",X"975962",X"973c79",
X"971f9f",X"9702d6",X"96e61d",X"96c975",X"96acdc",X"969054",X"9673dc",
X"965774",X"963b1d",X"961ed6",X"96029f",X"95e679",X"95ca63",X"95ae5d",
X"959268",X"957683",X"955aaf",X"953eeb",X"952337",X"950794",X"94ec02",
X"94d080",X"94b50e",X"9499ad",X"947e5d",X"94631d",X"9447ee",X"942ccf",
X"9411c1",X"93f6c4",X"93dbd7",X"93c0fb",X"93a630",X"938b75",X"9370cb",
X"935632",X"933baa",X"932132",X"9306cc",X"92ec76",X"92d230",X"92b7fc",
X"929dd9",X"9283c6",X"9269c4",X"924fd3",X"9235f3",X"921c24",X"920266",
X"91e8b9",X"91cf1d",X"91b592",X"919c18",X"9182af",X"916957",X"915010",
X"9136da",X"911db5",X"9104a1",X"90eb9f",X"90d2ad",X"90b9cd",X"90a0fe",
X"908840",X"906f93",X"9056f7",X"903e6d",X"9025f4",X"900d8c",X"8ff535",
X"8fdcf0",X"8fc4bc",X"8fac99",X"8f9488",X"8f7c88",X"8f6499",X"8f4cbb",
X"8f34ef",X"8f1d35",X"8f058c",X"8eedf4",X"8ed66d",X"8ebef8",X"8ea795",
X"8e9043",X"8e7903",X"8e61d4",X"8e4ab6",X"8e33aa",X"8e1cb0",X"8e05c7",
X"8deef0",X"8dd82a",X"8dc176",X"8daad4",X"8d9443",X"8d7dc4",X"8d6757",
X"8d50fb",X"8d3ab1",X"8d2478",X"8d0e52",X"8cf83d",X"8ce239",X"8ccc48",
X"8cb668",X"8ca09a",X"8c8ade",X"8c7534",X"8c5f9b",X"8c4a15",X"8c34a0",
X"8c1f3d",X"8c09ec",X"8bf4ad",X"8bdf7f",X"8bca64",X"8bb55a",X"8ba063",
X"8b8b7d",X"8b76a9",X"8b61e8",X"8b4d38",X"8b389a",X"8b240f",X"8b0f95",
X"8afb2d",X"8ae6d8",X"8ad294",X"8abe63",X"8aaa43",X"8a9636",X"8a823b",
X"8a6e52",X"8a5a7b",X"8a46b6",X"8a3303",X"8a1f63",X"8a0bd4",X"89f858",
X"89e4ee",X"89d197",X"89be51",X"89ab1e",X"8997fd",X"8984ee",X"8971f2",
X"895f08",X"894c30",X"89396a",X"8926b7",X"891416",X"890187",X"88ef0b",
X"88dca1",X"88ca4a",X"88b805",X"88a5d2",X"8893b2",X"8881a4",X"886fa8",
X"885dbf",X"884be9",X"883a24",X"882873",X"8816d4",X"880547",X"87f3cd",
X"87e265",X"87d110",X"87bfcd",X"87ae9d",X"879d80",X"878c75",X"877b7c",
X"876a97",X"8759c3",X"874903",X"873855",X"8727ba",X"871731",X"8706bb",
X"86f657",X"86e607",X"86d5c9",X"86c59d",X"86b584",X"86a57e",X"86958b",
X"8685ab",X"8675dd",X"866622",X"865679",X"8646e4",X"863761",X"8627f1",
X"861894",X"860949",X"85fa12",X"85eaed",X"85dbdb",X"85ccdc",X"85bdf0",
X"85af16",X"85a050",X"85919c",X"8582fb",X"85746d",X"8565f2",X"85578a",
X"854935",X"853af3",X"852cc3",X"851ea7",X"85109d",X"8502a7",X"84f4c3",
X"84e6f3",X"84d935",X"84cb8b",X"84bdf3",X"84b06e",X"84a2fd",X"84959e",
X"848853",X"847b1a",X"846df5",X"8460e3",X"8453e3",X"8446f7",X"843a1e",
X"842d58",X"8420a5",X"841405",X"840778",X"83faff",X"83ee98",X"83e245",
X"83d605",X"83c9d7",X"83bdbe",X"83b1b7",X"83a5c3",X"8399e3",X"838e16",
X"83825b",X"8376b5",X"836b21",X"835fa1",X"835433",X"8348d9",X"833d93",
X"83325f",X"83273f",X"831c32",X"831138",X"830652",X"82fb7e",X"82f0be",
X"82e612",X"82db78",X"82d0f2",X"82c680",X"82bc20",X"82b1d4",X"82a79b",
X"829d76",X"829364",X"828965",X"827f79",X"8275a1",X"826bdd",X"82622b",
X"82588d",X"824f03",X"82458b",X"823c27",X"8232d7",X"82299a",X"822070",
X"82175a",X"820e57",X"820568",X"81fc8c",X"81f3c3",X"81eb0e",X"81e26d",
X"81d9de",X"81d164",X"81c8fc",X"81c0a9",X"81b868",X"81b03b",X"81a822",
X"81a01c",X"819829",X"81904b",X"81887f",X"8180c7",X"817923",X"817192",
X"816a14",X"8162ab",X"815b54",X"815411",X"814ce2",X"8145c6",X"813ebe",
X"8137c9",X"8130e8",X"812a1b",X"812361",X"811cba",X"811627",X"810fa8",
X"81093c",X"8102e4",X"80fca0",X"80f66f",X"80f051",X"80ea48",X"80e451",
X"80de6f",X"80d8a0",X"80d2e4",X"80cd3d",X"80c7a9",X"80c228",X"80bcbb",
X"80b762",X"80b21c",X"80acea",X"80a7cc",X"80a2c1",X"809dca",X"8098e6",
X"809417",X"808f5b",X"808ab2",X"80861d",X"80819c",X"807d2e",X"8078d5",
X"80748e",X"80705c",X"806c3d",X"806832",X"80643a",X"806056",X"805c86",
X"8058ca",X"805521",X"80518c",X"804e0b",X"804a9d",X"804743",X"8043fc",
X"8040ca",X"803dab",X"803aa0",X"8037a8",X"8034c4",X"8031f4",X"802f38",
X"802c8f",X"8029fa",X"802779",X"80250b",X"8022b2",X"80206b",X"801e39",
X"801c1a",X"801a0f",X"801818",X"801635",X"801465",X"8012a9",X"801101",
X"800f6c",X"800deb",X"800c7e",X"800b25",X"8009df",X"8008ad",X"80078f",
X"800684",X"80058e",X"8004ab",X"8003db",X"800320",X"800278",X"8001e4",
X"800164",X"8000f7",X"80009e",X"800059",X"800028",X"80000a",X"800000",
X"80000a",X"800028",X"800059",X"80009e",X"8000f7",X"800164",X"8001e4",
X"800278",X"800320",X"8003db",X"8004ab",X"80058e",X"800684",X"80078f",
X"8008ad",X"8009df",X"800b25",X"800c7e",X"800deb",X"800f6c",X"801101",
X"8012a9",X"801465",X"801635",X"801818",X"801a0f",X"801c1a",X"801e39",
X"80206b",X"8022b2",X"80250b",X"802779",X"8029fa",X"802c8f",X"802f38",
X"8031f4",X"8034c4",X"8037a8",X"803aa0",X"803dab",X"8040ca",X"8043fc",
X"804743",X"804a9d",X"804e0b",X"80518c",X"805521",X"8058ca",X"805c86",
X"806056",X"80643a",X"806832",X"806c3d",X"80705c",X"80748e",X"8078d5",
X"807d2e",X"80819c",X"80861d",X"808ab2",X"808f5b",X"809417",X"8098e6",
X"809dca",X"80a2c1",X"80a7cc",X"80acea",X"80b21c",X"80b762",X"80bcbb",
X"80c228",X"80c7a9",X"80cd3d",X"80d2e4",X"80d8a0",X"80de6f",X"80e451",
X"80ea48",X"80f051",X"80f66f",X"80fca0",X"8102e4",X"81093c",X"810fa8",
X"811627",X"811cba",X"812361",X"812a1b",X"8130e8",X"8137c9",X"813ebe",
X"8145c6",X"814ce2",X"815411",X"815b54",X"8162ab",X"816a14",X"817192",
X"817923",X"8180c7",X"81887f",X"81904b",X"819829",X"81a01c",X"81a822",
X"81b03b",X"81b868",X"81c0a9",X"81c8fc",X"81d164",X"81d9de",X"81e26d",
X"81eb0e",X"81f3c3",X"81fc8c",X"820568",X"820e57",X"82175a",X"822070",
X"82299a",X"8232d7",X"823c27",X"82458b",X"824f03",X"82588d",X"82622b",
X"826bdd",X"8275a1",X"827f79",X"828965",X"829364",X"829d76",X"82a79b",
X"82b1d4",X"82bc20",X"82c680",X"82d0f2",X"82db78",X"82e612",X"82f0be",
X"82fb7e",X"830652",X"831138",X"831c32",X"83273f",X"83325f",X"833d93",
X"8348d9",X"835433",X"835fa1",X"836b21",X"8376b5",X"83825b",X"838e16",
X"8399e3",X"83a5c3",X"83b1b7",X"83bdbe",X"83c9d7",X"83d605",X"83e245",
X"83ee98",X"83faff",X"840778",X"841405",X"8420a5",X"842d58",X"843a1e",
X"8446f7",X"8453e3",X"8460e3",X"846df5",X"847b1a",X"848853",X"84959e",
X"84a2fd",X"84b06e",X"84bdf3",X"84cb8b",X"84d935",X"84e6f3",X"84f4c3",
X"8502a7",X"85109d",X"851ea7",X"852cc3",X"853af3",X"854935",X"85578a",
X"8565f2",X"85746d",X"8582fb",X"85919c",X"85a050",X"85af16",X"85bdf0",
X"85ccdc",X"85dbdb",X"85eaed",X"85fa12",X"860949",X"861894",X"8627f1",
X"863761",X"8646e4",X"865679",X"866622",X"8675dd",X"8685ab",X"86958b",
X"86a57e",X"86b584",X"86c59d",X"86d5c9",X"86e607",X"86f657",X"8706bb",
X"871731",X"8727ba",X"873855",X"874903",X"8759c3",X"876a97",X"877b7c",
X"878c75",X"879d80",X"87ae9d",X"87bfcd",X"87d110",X"87e265",X"87f3cd",
X"880547",X"8816d4",X"882873",X"883a24",X"884be9",X"885dbf",X"886fa8",
X"8881a4",X"8893b2",X"88a5d2",X"88b805",X"88ca4a",X"88dca1",X"88ef0b",
X"890187",X"891416",X"8926b7",X"89396a",X"894c30",X"895f08",X"8971f2",
X"8984ee",X"8997fd",X"89ab1e",X"89be51",X"89d197",X"89e4ee",X"89f858",
X"8a0bd4",X"8a1f63",X"8a3303",X"8a46b6",X"8a5a7b",X"8a6e52",X"8a823b",
X"8a9636",X"8aaa43",X"8abe63",X"8ad294",X"8ae6d8",X"8afb2d",X"8b0f95",
X"8b240f",X"8b389a",X"8b4d38",X"8b61e8",X"8b76a9",X"8b8b7d",X"8ba063",
X"8bb55a",X"8bca64",X"8bdf7f",X"8bf4ad",X"8c09ec",X"8c1f3d",X"8c34a0",
X"8c4a15",X"8c5f9b",X"8c7534",X"8c8ade",X"8ca09a",X"8cb668",X"8ccc48",
X"8ce239",X"8cf83d",X"8d0e52",X"8d2478",X"8d3ab1",X"8d50fb",X"8d6757",
X"8d7dc4",X"8d9443",X"8daad4",X"8dc176",X"8dd82a",X"8deef0",X"8e05c7",
X"8e1cb0",X"8e33aa",X"8e4ab6",X"8e61d4",X"8e7903",X"8e9043",X"8ea795",
X"8ebef8",X"8ed66d",X"8eedf4",X"8f058c",X"8f1d35",X"8f34ef",X"8f4cbb",
X"8f6499",X"8f7c88",X"8f9488",X"8fac99",X"8fc4bc",X"8fdcf0",X"8ff535",
X"900d8c",X"9025f4",X"903e6d",X"9056f7",X"906f93",X"908840",X"90a0fe",
X"90b9cd",X"90d2ad",X"90eb9f",X"9104a1",X"911db5",X"9136da",X"915010",
X"916957",X"9182af",X"919c18",X"91b592",X"91cf1d",X"91e8b9",X"920266",
X"921c24",X"9235f3",X"924fd3",X"9269c4",X"9283c6",X"929dd9",X"92b7fc",
X"92d230",X"92ec76",X"9306cc",X"932132",X"933baa",X"935632",X"9370cb",
X"938b75",X"93a630",X"93c0fb",X"93dbd7",X"93f6c4",X"9411c1",X"942ccf",
X"9447ee",X"94631d",X"947e5d",X"9499ad",X"94b50e",X"94d080",X"94ec02",
X"950794",X"952337",X"953eeb",X"955aaf",X"957683",X"959268",X"95ae5d",
X"95ca63",X"95e679",X"96029f",X"961ed6",X"963b1d",X"965774",X"9673dc",
X"969054",X"96acdc",X"96c975",X"96e61d",X"9702d6",X"971f9f",X"973c79",
X"975962",X"97765c",X"979365",X"97b07f",X"97cda9",X"97eae3",X"98082d",
X"982587",X"9842f1",X"98606b",X"987df5",X"989b8f",X"98b939",X"98d6f2",
X"98f4bc",X"991296",X"99307f",X"994e79",X"996c82",X"998a9b",X"99a8c4",
X"99c6fc",X"99e545",X"9a039d",X"9a2205",X"9a407c",X"9a5f03",X"9a7d9a",
X"9a9c41",X"9abaf7",X"9ad9bd",X"9af892",X"9b1777",X"9b366c",X"9b5570",
X"9b7484",X"9b93a7",X"9bb2d9",X"9bd21b",X"9bf16d",X"9c10ce",X"9c303e",
X"9c4fbe",X"9c6f4d",X"9c8eec",X"9cae9a",X"9cce57",X"9cee23",X"9d0dff",
X"9d2dea",X"9d4de4",X"9d6ded",X"9d8e06",X"9dae2e",X"9dce65",X"9deeab",
X"9e0f00",X"9e2f65",X"9e4fd8",X"9e705b",X"9e90ec",X"9eb18d",X"9ed23c",
X"9ef2fb",X"9f13c8",X"9f34a5",X"9f5590",X"9f768a",X"9f9794",X"9fb8ac",
X"9fd9d3",X"9ffb08",X"a01c4d",X"a03da0",X"a05f02",X"a08073",X"a0a1f3",
X"a0c381",X"a0e51e",X"a106ca",X"a12884",X"a14a4d",X"a16c24",X"a18e0a",
X"a1afff",X"a1d202",X"a1f414",X"a21634",X"a23863",X"a25aa0",X"a27cec",
X"a29f46",X"a2c1ae",X"a2e425",X"a306aa",X"a3293e",X"a34be0",X"a36e90",
X"a3914e",X"a3b41b",X"a3d6f6",X"a3f9df",X"a41cd6",X"a43fdc",X"a462ef",
X"a48611",X"a4a941",X"a4cc7f",X"a4efcb",X"a51325",X"a5368d",X"a55a03",
X"a57d87",X"a5a119",X"a5c4b9",X"a5e867",X"a60c22",X"a62fec",X"a653c4",
X"a677a9",X"a69b9c",X"a6bf9d",X"a6e3ab",X"a707c8",X"a72bf2",X"a7502a",
X"a7746f",X"a798c2",X"a7bd23",X"a7e192",X"a8060e",X"a82a97",X"a84f2e",
X"a873d3",X"a89885",X"a8bd44",X"a8e212",X"a906ec",X"a92bd4",X"a950c9",
X"a975cc",X"a99adc",X"a9bff9",X"a9e524",X"aa0a5c",X"aa2fa1",X"aa54f3",
X"aa7a53",X"aa9fc0",X"aac53a",X"aaeac1",X"ab1055",X"ab35f6",X"ab5ba5",
X"ab8160",X"aba729",X"abccfe",X"abf2e0",X"ac18d0",X"ac3ecc",X"ac64d6",
X"ac8aec",X"acb10f",X"acd73f",X"acfd7b",X"ad23c5",X"ad4a1b",X"ad707e",
X"ad96ee",X"adbd6b",X"ade3f4",X"ae0a8a",X"ae312c",X"ae57db",X"ae7e97",
X"aea55f",X"aecc34",X"aef315",X"af1a03",X"af40fd",X"af6804",X"af8f17",
X"afb637",X"afdd63",X"b0049b",X"b02be0",X"b05331",X"b07a8e",X"b0a1f8",
X"b0c96d",X"b0f0ef",X"b1187e",X"b14018",X"b167be",X"b18f71",X"b1b730",
X"b1defa",X"b206d1",X"b22eb4",X"b256a3",X"b27e9e",X"b2a6a5",X"b2ceb7",
X"b2f6d6",X"b31f00",X"b34737",X"b36f79",X"b397c7",X"b3c021",X"b3e886",
X"b410f7",X"b43974",X"b461fd",X"b48a91",X"b4b331",X"b4dbdd",X"b50494",
X"b52d57",X"b55625",X"b57eff",X"b5a7e4",X"b5d0d5",X"b5f9d1",X"b622d8",
X"b64beb",X"b6750a",X"b69e33",X"b6c768",X"b6f0a9",X"b719f4",X"b7434b",
X"b76cad",X"b7961a",X"b7bf92",X"b7e916",X"b812a5",X"b83c3e",X"b865e3",
X"b88f93",X"b8b94e",X"b8e314",X"b90ce4",X"b936c0",X"b960a7",X"b98a98",
X"b9b495",X"b9de9c",X"ba08ae",X"ba32cb",X"ba5cf3",X"ba8725",X"bab162",
X"badbaa",X"bb05fc",X"bb3059",X"bb5ac1",X"bb8533",X"bbafb0",X"bbda37",
X"bc04c9",X"bc2f66",X"bc5a0c",X"bc84be",X"bcaf79",X"bcda3f",X"bd0510",
X"bd2fea",X"bd5acf",X"bd85bf",X"bdb0b8",X"bddbbc",X"be06ca",X"be31e2",
X"be5d04",X"be8831",X"beb367",X"bedea8",X"bf09f3",X"bf3547",X"bf60a6",
X"bf8c0e",X"bfb781",X"bfe2fd",X"c00e84",X"c03a14",X"c065ae",X"c09152",
X"c0bcff",X"c0e8b7",X"c11478",X"c14043",X"c16c17",X"c197f5",X"c1c3dd",
X"c1efce",X"c21bc9",X"c247ce",X"c273dc",X"c29ff3",X"c2cc14",X"c2f83f",
X"c32472",X"c350b0",X"c37cf6",X"c3a946",X"c3d59f",X"c40202",X"c42e6d",
X"c45ae2",X"c48760",X"c4b3e8",X"c4e078",X"c50d12",X"c539b4",X"c56660",
X"c59315",X"c5bfd3",X"c5ec99",X"c61969",X"c64642",X"c67323",X"c6a00e",
X"c6cd01",X"c6f9fd",X"c72702",X"c75410",X"c78126",X"c7ae45",X"c7db6d",
X"c8089d",X"c835d6",X"c86318",X"c89062",X"c8bdb5",X"c8eb10",X"c91874",
X"c945e0",X"c97355",X"c9a0d2",X"c9ce58",X"c9fbe6",X"ca297c",X"ca571a",
X"ca84c1",X"cab270",X"cae027",X"cb0de7",X"cb3bae",X"cb697e",X"cb9756",
X"cbc536",X"cbf31e",X"cc210e",X"cc4f06",X"cc7d06",X"ccab0e",X"ccd91e",
X"cd0735",X"cd3555",X"cd637c",X"cd91ac",X"cdbfe3",X"cdee21",X"ce1c68",
X"ce4ab6",X"ce790c",X"cea769",X"ced5cf",X"cf043b",X"cf32af",X"cf612b",
X"cf8fae",X"cfbe39",X"cfeccb",X"d01b65",X"d04a06",X"d078ae",X"d0a75e",
X"d0d615",X"d104d3",X"d13398",X"d16265",X"d19139",X"d1c014",X"d1eef6",
X"d21ddf",X"d24cd0",X"d27bc7",X"d2aac6",X"d2d9cb",X"d308d7",X"d337eb",
X"d36705",X"d39626",X"d3c54e",X"d3f47d",X"d423b2",X"d452ee",X"d48231",
X"d4b17b",X"d4e0cc",X"d51023",X"d53f80",X"d56ee5",X"d59e4f",X"d5cdc1",
X"d5fd39",X"d62cb7",X"d65c3c",X"d68bc7",X"d6bb59",X"d6eaf1",X"d71a8f",
X"d74a34",X"d779df",X"d7a990",X"d7d947",X"d80905",X"d838c9",X"d86893",
X"d89863",X"d8c839",X"d8f815",X"d927f7",X"d957df",X"d987cd",X"d9b7c1",
X"d9e7bb",X"da17bb",X"da47c0",X"da77cc",X"daa7dd",X"dad7f4",X"db0811",
X"db3833",X"db685b",X"db9889",X"dbc8bd",X"dbf8f5",X"dc2934",X"dc5978",
X"dc89c2",X"dcba11",X"dcea65",X"dd1abf",X"dd4b1e",X"dd7b83",X"ddabed",
X"dddc5c",X"de0cd0",X"de3d4a",X"de6dc9",X"de9e4d",X"deced6",X"deff64",
X"df2ff8",X"df6090",X"df912e",X"dfc1d0",X"dff278",X"e02324",X"e053d6",
X"e0848c",X"e0b547",X"e0e607",X"e116cc",X"e14795",X"e17863",X"e1a936",
X"e1da0e",X"e20aea",X"e23bcb",X"e26cb1",X"e29d9b",X"e2ce89",X"e2ff7c",
X"e33074",X"e36170",X"e39270",X"e3c375",X"e3f47e",X"e4258c",X"e4569d",
X"e487b3",X"e4b8ce",X"e4e9ec",X"e51b0f",X"e54c35",X"e57d60",X"e5ae8f",
X"e5dfc2",X"e610f9",X"e64235",X"e67374",X"e6a4b7",X"e6d5fd",X"e70748",
X"e73897",X"e769e9",X"e79b40",X"e7cc9a",X"e7fdf7",X"e82f59",X"e860be",
X"e89227",X"e8c393",X"e8f503",X"e92676",X"e957ed",X"e98968",X"e9bae6",
X"e9ec67",X"ea1dec",X"ea4f74",X"ea8100",X"eab28f",X"eae421",X"eb15b6",
X"eb474f",X"eb78eb",X"ebaa8a",X"ebdc2c",X"ec0dd1",X"ec3f79",X"ec7125",
X"eca2d3",X"ecd485",X"ed0639",X"ed37f0",X"ed69aa",X"ed9b67",X"edcd27",
X"edfeea",X"ee30af",X"ee6277",X"ee9442",X"eec610",X"eef7e0",X"ef29b3",
X"ef5b88",X"ef8d60",X"efbf3b",X"eff118",X"f022f7",X"f054d9",X"f086be",
X"f0b8a5",X"f0ea8e",X"f11c79",X"f14e67",X"f18057",X"f1b249",X"f1e43e",
X"f21634",X"f2482d",X"f27a28",X"f2ac25",X"f2de24",X"f31025",X"f34228",
X"f3742d",X"f3a634",X"f3d83d",X"f40a48",X"f43c54",X"f46e63",X"f4a073",
X"f4d285",X"f50498",X"f536ae",X"f568c5",X"f59ade",X"f5ccf8",X"f5ff14",
X"f63131",X"f66350",X"f69570",X"f6c792",X"f6f9b5",X"f72bda",X"f75e00",
X"f79027",X"f7c250",X"f7f47a",X"f826a5",X"f858d1",X"f88aff",X"f8bd2d",
X"f8ef5d",X"f9218e",X"f953c0",X"f985f3",X"f9b827",X"f9ea5c",X"fa1c92",
X"fa4ec9",X"fa8100",X"fab339",X"fae572",X"fb17ac",X"fb49e7",X"fb7c23",
X"fbae5f",X"fbe09c",X"fc12da",X"fc4518",X"fc7757",X"fca996",X"fcdbd6",
X"fd0e16",X"fd4057",X"fd7298",X"fda4da",X"fdd71c",X"fe095e",X"fe3ba1",
X"fe6de3",X"fea026",X"fed26a",X"ff04ad",X"ff36f1",X"ff6935",X"ff9b79",
X"ffcdbd"
);

begin

rom_select: process (clk)
begin
	if clk'event and clk = '1' then
		if en = '1' then
			sin_out <= sin_ROM(conv_integer(addr));
		end if;
	end if;
end process rom_select;
end rtl;